module fifo #(
    parameter DATA_WIDTH = 8,
    parameter DEPTH 	= 16
) (
    input wire i_Clock,
    input wire i_reset,
    input wire wr_en,
    input wire rd_en,
    input wire [DATA_WIDTH-1:0] data_in,
    output wire [DATA_WIDTH-1:0] data_out,
    output wire full,
    output wire empty
);

	 reg [DATA_WIDTH-1:0] mem [0:DEPTH-1];
	 reg [4:0] rd_ptr, wr_ptr;
	 reg [4:0] count;

	 assign data_out = mem[rd_ptr];
	 assign full  = (count == DEPTH);
	 assign empty = (count == 0);

always @(posedge i_Clock or negedge i_reset) begin
    if (~i_reset) begin
        rd_ptr <= 0;
        wr_ptr <= 0;
        count <= 0;
    end else begin
        if (wr_en & ~full) begin
            mem[wr_ptr] <= data_in;
            wr_ptr <= wr_ptr + 1;
            count <= count + 1;
        end
        if (rd_en & ~empty) begin
            rd_ptr <= rd_ptr + 1;
            count <= count - 1;
        end
    end
end

endmodule
